  ***project_cmos(created by dharmendra)

.subckt invertor_ckt 1 2 3
.model nmod nmos level=54 version=4.7
.model pmod pmos level=54 version=4.7
M1 3 1 0 0 nmod w=100u l=10u
M2 3 1 2 2 pmod w=100u l=10u
.ends

.subckt NAND_CKT 1 2 3 4 
.model nmod nmos level=54 version=4.7
.model pmod pmos level=54 version=4.7
M1 5 1 0 0 nmod w=100u l=10u
M2 4 2 5 5 nmod w=100u l=10u
M3 4 2 3 3 pmod w=100u l=10u
M4 4 1 3 3 pmod w=100l l=10u
.ends

.subbckt XOR_CKT 11 12 16
Xfirst_nand 11 12 2 13 NAND_CKT
Xsecond_nand 12 13 2 14 NAND_CKT
Xthird_nand 11 13 2 15 NAND_CKT
Xfourth_nand 14 15 2 16 NAND_CKT
.ends 

.subckt MUX_CKT 11 12 13 17
Xfirst_nand 11 13 2 15 NAND_CKT
Xinvert 13 2 14 invertor_ckt
Xsecond_nand 12 14 2 16 NAND_CKT
Xthird_nand 15 16 2 17 NAND_CKT
.ends

Va 21 0 dc 0v 
Vb 22 0 dc 0v 
Vc 24 0 dc 0v 
Vd 25 0 pulse(0 5 0 0 0 10m 20m)
Ve 29 0 dc 0v
Vdd 2 0 dc 5v

Xxor_1 21 22 23 XOR_CKT
Xxor_2 24 25 27 XOR_CKT
Xmux_1 21 24 23 26 MUX_CKT
Xxor_3 23 27 28 XOR_CKT
Xmux_2 25 28 29 31 MUX_CKT
Xxor_4 28 29 30 XOR_CKT

.tran 0.1m 100m 
.control
run
plot V(31)
plot V(30)
plot V(26)
.endc
.end


